/*
==============================================
* SAR Assertions and Coverage
    To be bound with SAR Top.
*   Date: 4/25/24
==============================================
*/

import tst_config_pkg::*;
module sar_ac (
    dbe_if.dut dbe,
    afe_if afe
);


endmodule
